VERSION 5.8 ;
BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

MACRO UART
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  SIZE 48.712 BY 47.8 ;
  SYMMETRY X Y ;
  PIN RST
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 22.428 0 22.484 0.286 ;
    END
  END RST
  PIN TX_CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M4 ;
        RECT 20.908 0 20.964 0.286 ;
    END
  END TX_CLK
  PIN RX_CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M3 ;
        RECT 0 24.252 0.286 24.308 ;
    END
  END RX_CLK
  PIN RX_IN_S
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 30.332 47.514 30.388 47.8 ;
    END
  END RX_IN_S
  PIN RX_OUT_P[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 48.426 35.196 48.712 35.252 ;
    END
  END RX_OUT_P[7]
  PIN RX_OUT_P[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 48.426 37.628 48.712 37.684 ;
    END
  END RX_OUT_P[6]
  PIN RX_OUT_P[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 48.426 35.5 48.712 35.556 ;
    END
  END RX_OUT_P[5]
  PIN RX_OUT_P[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 48.426 39.756 48.712 39.812 ;
    END
  END RX_OUT_P[4]
  PIN RX_OUT_P[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 41.58 47.514 41.636 47.8 ;
    END
  END RX_OUT_P[3]
  PIN RX_OUT_P[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 38.844 47.514 38.9 47.8 ;
    END
  END RX_OUT_P[2]
  PIN RX_OUT_P[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 36.716 47.514 36.772 47.8 ;
    END
  END RX_OUT_P[1]
  PIN RX_OUT_P[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 34.588 47.514 34.644 47.8 ;
    END
  END RX_OUT_P[0]
  PIN RX_OUT_V
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 48.426 28.812 48.712 28.868 ;
    END
  END RX_OUT_V
  PIN TX_IN_P[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 29.724 0 29.78 0.286 ;
    END
  END TX_IN_P[7]
  PIN TX_IN_P[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 27.292 0 27.348 0.286 ;
    END
  END TX_IN_P[6]
  PIN TX_IN_P[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 27.9 0 27.956 0.286 ;
    END
  END TX_IN_P[5]
  PIN TX_IN_P[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 25.772 0 25.828 0.286 ;
    END
  END TX_IN_P[4]
  PIN TX_IN_P[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 32.156 0 32.212 0.286 ;
    END
  END TX_IN_P[3]
  PIN TX_IN_P[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 48.426 18.172 48.712 18.228 ;
    END
  END TX_IN_P[2]
  PIN TX_IN_P[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 30.028 0 30.084 0.286 ;
    END
  END TX_IN_P[1]
  PIN TX_IN_P[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16.652 0 16.708 0.286 ;
    END
  END TX_IN_P[0]
  PIN TX_IN_V
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 32.764 0 32.82 0.286 ;
    END
  END TX_IN_V
  PIN TX_OUT_S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 48.426 16.044 48.712 16.1 ;
    END
  END TX_OUT_S
  PIN TX_OUT_V
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 34.892 0 34.948 0.286 ;
    END
  END TX_OUT_V
  PIN Prescale[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0 21.82 0.286 21.876 ;
    END
  END Prescale[5]
  PIN Prescale[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0 14.828 0.286 14.884 ;
    END
  END Prescale[4]
  PIN Prescale[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0 26.38 0.286 26.436 ;
    END
  END Prescale[3]
  PIN Prescale[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0 21.516 0.286 21.572 ;
    END
  END Prescale[2]
  PIN Prescale[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0 28.508 0.286 28.564 ;
    END
  END Prescale[1]
  PIN Prescale[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0 18.78 0.286 18.836 ;
    END
  END Prescale[0]
  PIN parity_enable
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 48.426 19.388 48.712 19.444 ;
    END
  END parity_enable
  PIN parity_type
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 48.426 21.82 48.712 21.876 ;
    END
  END parity_type
  PIN parity_error
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 48.426 30.94 48.712 30.996 ;
    END
  END parity_error
  PIN framing_error
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 48.426 26.684 48.712 26.74 ;
    END
  END framing_error
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13.612 47.514 13.668 47.8 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 24.556 47.514 24.612 47.8 ;
    END
  END SE
  PIN SO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 48.426 23.948 48.712 24.004 ;
    END
  END SO
  PIN scan_clk
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M4 ;
        RECT 18.78 0 18.836 0.286 ;
    END
  END scan_clk
  PIN scan_rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 23.036 0 23.092 0.286 ;
    END
  END scan_rst
  PIN test_mode
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 24.86 0 24.916 0.286 ;
    END
  END test_mode
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
  END VSS
  OBS
    LAYER M6 ;
      RECT 23.184 0.7 24.16 1.005 ;
      RECT 25.616 0.7 26.592 1.005 ;
      RECT 28.048 0.7 29.024 1.005 ;
      RECT 30.48 0.7 31.456 1.005 ;
      RECT 0.7 0.986 48.012 47.1 ;
      RECT 0.7 0.7 21.728 3.705 ;
      RECT 32.912 0.7 48.012 3.705 ;
    LAYER M4 ;
      RECT 35.344 46.795 36.016 47.1 ;
      RECT 37.472 46.795 38.144 47.1 ;
      RECT 39.6 46.795 40.88 47.1 ;
      RECT 17.408 0.7 18.08 1.005 ;
      RECT 19.536 0.7 20.208 1.005 ;
      RECT 21.664 0.7 22.336 1.005 ;
      RECT 23.792 0.7 25.072 1.005 ;
      RECT 26.528 0.7 27.2 1.005 ;
      RECT 28.656 0.7 29.328 1.005 ;
      RECT 30.784 0.7 32.064 1.005 ;
      RECT 33.52 0.7 34.192 1.005 ;
      RECT 31.088 45.595 33.888 47.1 ;
      RECT 0.7 44.095 12.912 47.1 ;
      RECT 14.368 44.095 23.856 47.1 ;
      RECT 25.312 44.095 29.632 47.1 ;
      RECT 42.336 44.095 48.012 47.1 ;
      RECT 0.7 0.986 48.012 46.814 ;
      RECT 0.7 0.7 15.952 3.705 ;
      RECT 35.648 0.7 48.012 3.705 ;
      POLYGON 48.012 47.1 48.012 0.7 35.648 0.7 35.648 0.986 34.192 0.986 34.192 0.7 33.52 0.7 33.52 0.986 32.064 0.986 32.064 0.7 30.784 0.7 30.784 0.986 29.328 0.986 29.328 0.7 28.656 0.7 28.656 0.986 27.2 0.986 27.2 0.7 26.528 0.7 26.528 0.986 25.072 0.986 25.072 0.7 24.308 0.7 24.308 0.623 24.31 0.623 24.31 0.513 24.25 0.513 24.25 0.623 24.252 0.623 24.252 0.7 23.792 0.7 23.792 0.986 22.336 0.986 22.336 0.7 21.664 0.7 21.664 0.986 20.208 0.986 20.208 0.7 19.536 0.7 19.536 0.986 18.08 0.986 18.08 0.7 17.408 0.7 17.408 0.986 15.952 0.986 15.952 0.7 0.7 0.7 0.7 47.1 12.912 47.1 12.912 46.814 14.368 46.814 14.368 47.1 23.856 47.1 23.856 46.814 25.312 46.814 25.312 47.1 29.632 47.1 29.632 46.814 31.088 46.814 31.088 47.1 33.888 47.1 33.888 46.814 35.344 46.814 35.344 47.1 36.016 47.1 36.016 46.814 37.472 46.814 37.472 47.1 38.144 47.1 38.144 46.814 39.6 46.814 39.6 47.1 40.88 47.1 40.88 46.814 42.336 46.814 42.336 47.1 ;
      POLYGON 48.63 19.471 48.63 19.361 48.628 19.361 48.628 18.863 48.63 18.863 48.63 18.753 48.57 18.753 48.57 18.863 48.572 18.863 48.572 19.361 48.57 19.361 48.57 19.471 ;
    LAYER M3 ;
      RECT 47.707 38.384 48.012 39.056 ;
      RECT 47.707 36.256 48.012 36.928 ;
      RECT 47.707 29.568 48.012 30.24 ;
      RECT 47.707 27.44 48.012 28.112 ;
      RECT 0.7 27.136 1.005 27.808 ;
      RECT 47.707 24.704 48.012 25.984 ;
      RECT 0.7 25.008 1.005 25.68 ;
      RECT 0.7 22.272 1.005 23.552 ;
      RECT 47.707 22.576 48.012 23.248 ;
      RECT 0.7 19.536 1.005 20.816 ;
      RECT 47.707 16.8 48.012 17.472 ;
      RECT 46.507 18.928 48.012 21.12 ;
      RECT 0.7 15.584 2.205 18.08 ;
      RECT 0.7 40.512 48.012 47.1 ;
      RECT 0.7 34.8 47.726 40.512 ;
      RECT 0.7 31.696 48.012 34.8 ;
      RECT 0.7 29.264 47.726 32.269 ;
      RECT 0.986 15.344 47.726 29.264 ;
      RECT 0.986 14.128 47.726 17.133 ;
      RECT 45.007 12.339 48.012 15.344 ;
      RECT 0.7 0.7 48.012 14.128 ;
      POLYGON 48.012 47.1 48.012 40.512 47.726 40.512 47.726 39.056 48.012 39.056 48.012 38.384 47.726 38.384 47.726 36.928 48.012 36.928 48.012 36.256 47.726 36.256 47.726 34.8 48.012 34.8 48.012 31.696 47.726 31.696 47.726 30.24 48.012 30.24 48.012 29.568 47.726 29.568 47.726 28.112 48.012 28.112 48.012 27.44 47.726 27.44 47.726 25.984 48.012 25.984 48.012 24.704 47.726 24.704 47.726 23.248 48.012 23.248 48.012 22.576 47.726 22.576 47.726 21.12 48.012 21.12 48.012 18.928 47.726 18.928 47.726 18.836 48.545 18.836 48.545 18.838 48.655 18.838 48.655 18.778 48.545 18.778 48.545 18.78 47.726 18.78 47.726 17.472 48.012 17.472 48.012 16.8 47.726 16.8 47.726 15.344 48.012 15.344 48.012 0.7 0.7 0.7 0.7 14.128 0.986 14.128 0.986 15.584 0.7 15.584 0.7 18.08 0.986 18.08 0.986 19.536 0.7 19.536 0.7 20.816 0.986 20.816 0.986 22.272 0.7 22.272 0.7 23.552 0.986 23.552 0.986 25.008 0.7 25.008 0.7 25.68 0.986 25.68 0.986 27.136 0.7 27.136 0.7 27.808 0.986 27.808 0.986 29.264 0.7 29.264 0.7 47.1 ;
      POLYGON 27.983 0.598 27.983 0.538 27.873 0.538 27.873 0.54 22.967 0.54 22.967 0.538 22.857 0.538 22.857 0.598 22.967 0.598 22.967 0.596 27.873 0.596 27.873 0.598 ;
    LAYER M5 ;
      RECT 0.7 35.952 48.012 47.1 ;
      RECT 0.7 32.947 47.726 37.501 ;
      RECT 0.7 22.576 48.012 34.496 ;
      RECT 0.986 20.144 48.012 24.125 ;
      RECT 0.986 21.071 48.012 22.576 ;
      RECT 0.7 18.115 3.705 21.12 ;
      RECT 3.705 20.144 48.012 23.149 ;
      RECT 0.986 18.688 47.726 21.693 ;
      RECT 0.7 18.115 3.705 21.12 ;
      RECT 0.7 0.7 48.012 18.688 ;
      POLYGON 48.012 47.1 48.012 35.952 47.726 35.952 47.726 34.496 48.012 34.496 48.012 20.144 47.726 20.144 47.726 18.688 48.012 18.688 48.012 0.7 0.7 0.7 0.7 21.12 0.986 21.12 0.986 22.576 0.7 22.576 0.7 47.1 ;
      POLYGON 27.375 0.598 27.375 0.538 27.265 0.538 27.265 0.54 24.335 0.54 24.335 0.538 24.225 0.538 24.225 0.598 24.335 0.598 24.335 0.596 27.265 0.596 27.265 0.598 ;
    LAYER NWELL ;
      RECT 0.23 0.23 48.482 47.57 ;
    LAYER PO ;
      RECT 0.122 0.122 48.59 47.678 ;
    LAYER M1 ;
      RECT 0.6 0.6 48.112 47.2 ;
    LAYER M2 ;
      RECT 0.7 0.7 48.012 47.1 ;
      POLYGON 48.012 47.1 48.012 0.7 22.94 0.7 22.94 0.623 22.942 0.623 22.942 0.513 22.882 0.513 22.882 0.623 22.884 0.623 22.884 0.7 0.7 0.7 0.7 47.1 ;
    LAYER VIA2 ;
      RECT 22.887 0.543 22.937 0.593 ;
    LAYER VIA3 ;
      RECT 0.847 24.255 0.897 24.305 ;
      RECT 48.575 18.783 48.625 18.833 ;
      RECT 27.903 0.543 27.953 0.593 ;
    LAYER VIA4 ;
      RECT 48.575 19.391 48.625 19.441 ;
      RECT 24.255 0.543 24.305 0.593 ;
    LAYER VIA5 ;
      RECT 27.295 0.543 27.345 0.593 ;
    LAYER M7 ;
      RECT 0.7 0.7 48.012 47.1 ;
    LAYER M8 ;
      RECT 0.7 0.7 48.012 47.1 ;
    LAYER M9 ;
      RECT 0.5 0.5 48.212 47.3 ;
    LAYER MRDL ;
      RECT 2 2 46.712 45.8 ;
    LAYER OVERLAP ;
      POLYGON 0 0 0 47.8 48.712 47.8 48.712 0 ;
  END
END UART

END LIBRARY
