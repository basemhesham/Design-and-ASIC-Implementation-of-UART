VERSION 5.8 ;
BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

MACRO UART
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  SIZE 56.056 BY 55.144 ;
  SYMMETRY X Y ;
  PIN RST
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 24.732 0 24.788 0.286 ;
    END
  END RST
  PIN TX_CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M6 ;
        RECT 25.644 0 25.7 0.286 ;
    END
  END TX_CLK
  PIN RX_CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M3 ;
        RECT 0 27.164 0.286 27.22 ;
    END
  END RX_CLK
  PIN RX_IN_S
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 33.244 54.858 33.3 55.144 ;
    END
  END RX_IN_S
  PIN RX_OUT_P[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 55.77 45.708 56.056 45.764 ;
    END
  END RX_OUT_P[7]
  PIN RX_OUT_P[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 55.77 39.02 56.056 39.076 ;
    END
  END RX_OUT_P[6]
  PIN RX_OUT_P[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 55.77 41.148 56.056 41.204 ;
    END
  END RX_OUT_P[5]
  PIN RX_OUT_P[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 55.77 43.58 56.056 43.636 ;
    END
  END RX_OUT_P[4]
  PIN RX_OUT_P[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 46.924 54.858 46.98 55.144 ;
    END
  END RX_OUT_P[3]
  PIN RX_OUT_P[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 43.276 54.858 43.332 55.144 ;
    END
  END RX_OUT_P[2]
  PIN RX_OUT_P[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 41.148 54.858 41.204 55.144 ;
    END
  END RX_OUT_P[1]
  PIN RX_OUT_P[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 39.02 54.858 39.076 55.144 ;
    END
  END RX_OUT_P[0]
  PIN RX_OUT_V
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 55.77 34.156 56.056 34.212 ;
    END
  END RX_OUT_V
  PIN TX_IN_P[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 34.764 0 34.82 0.286 ;
    END
  END TX_IN_P[7]
  PIN TX_IN_P[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 31.724 0 31.78 0.286 ;
    END
  END TX_IN_P[6]
  PIN TX_IN_P[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 31.116 0 31.172 0.286 ;
    END
  END TX_IN_P[5]
  PIN TX_IN_P[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 20.476 0 20.532 0.286 ;
    END
  END TX_IN_P[4]
  PIN TX_IN_P[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 28.076 0 28.132 0.286 ;
    END
  END TX_IN_P[3]
  PIN TX_IN_P[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 55.77 21.084 56.056 21.14 ;
    END
  END TX_IN_P[2]
  PIN TX_IN_P[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 33.244 0 33.3 0.286 ;
    END
  END TX_IN_P[1]
  PIN TX_IN_P[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 35.372 0 35.428 0.286 ;
    END
  END TX_IN_P[0]
  PIN TX_IN_V
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 41.148 0 41.204 0.286 ;
    END
  END TX_IN_V
  PIN TX_OUT_S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 55.77 23.212 56.056 23.268 ;
    END
  END TX_OUT_S
  PIN TX_OUT_V
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 39.02 0 39.076 0.286 ;
    END
  END TX_OUT_V
  PIN Prescale[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0 23.516 0.286 23.572 ;
    END
  END Prescale[5]
  PIN Prescale[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0 20.172 0.286 20.228 ;
    END
  END Prescale[4]
  PIN Prescale[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0 31.42 0.286 31.476 ;
    END
  END Prescale[3]
  PIN Prescale[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0 26.86 0.286 26.916 ;
    END
  END Prescale[2]
  PIN Prescale[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0 33.548 0.286 33.604 ;
    END
  END Prescale[1]
  PIN Prescale[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0 29.292 0.286 29.348 ;
    END
  END Prescale[0]
  PIN parity_enable
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 55.77 18.956 56.056 19.012 ;
    END
  END parity_enable
  PIN parity_type
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 55.77 26.556 56.056 26.612 ;
    END
  END parity_type
  PIN parity_error
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 55.77 32.028 56.056 32.084 ;
    END
  END parity_error
  PIN framing_error
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 55.77 36.284 56.056 36.34 ;
    END
  END framing_error
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16.22 54.858 16.276 55.144 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 26.556 54.858 26.612 55.144 ;
    END
  END SE
  PIN SO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 55.77 29.292 56.056 29.348 ;
    END
  END SO
  PIN scan_clk
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M4 ;
        RECT 28.988 0 29.044 0.286 ;
    END
  END scan_clk
  PIN scan_rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 26.86 0 26.916 0.286 ;
    END
  END scan_rst
  PIN test_mode
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 22.604 0 22.66 0.286 ;
    END
  END test_mode
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER M9 ;
        RECT 0 3 1 4 ;
        RECT 55.056 3 56.056 4 ;
        RECT 0 51.144 1 52.144 ;
        RECT 55.056 51.144 56.056 52.144 ;
      LAYER M8 ;
        RECT 3 0 4 1 ;
        RECT 52.056 0 53.056 1 ;
        RECT 3 54.144 4 55.144 ;
        RECT 52.056 54.144 53.056 55.144 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER M9 ;
        RECT 0 1.6 1 2.6 ;
        RECT 55.056 1.6 56.056 2.6 ;
        RECT 0 52.544 1 53.544 ;
        RECT 55.056 52.544 56.056 53.544 ;
      LAYER M8 ;
        RECT 1.6 0 2.6 1 ;
        RECT 53.456 0 54.456 1 ;
        RECT 1.6 54.144 2.6 55.144 ;
        RECT 53.456 54.144 54.456 55.144 ;
    END
  END VSS
  OBS
    LAYER M4 ;
      RECT 39.776 54.139 40.448 54.444 ;
      RECT 41.904 54.139 42.576 54.444 ;
      RECT 21.232 0.7 21.904 1.005 ;
      RECT 23.36 0.7 24.032 1.005 ;
      RECT 25.488 0.7 26.16 1.005 ;
      RECT 27.616 0.7 28.288 1.005 ;
      RECT 29.744 0.7 30.416 1.005 ;
      RECT 31.872 0.7 32.544 1.005 ;
      RECT 34 0.7 34.672 1.005 ;
      RECT 39.776 0.7 40.448 1.005 ;
      RECT 44.032 52.939 46.224 54.444 ;
      RECT 36.128 0.7 38.32 2.205 ;
      RECT 0.7 51.439 15.52 54.444 ;
      RECT 16.976 51.439 25.856 54.444 ;
      RECT 27.312 51.439 32.544 54.444 ;
      RECT 34 51.439 38.32 54.444 ;
      RECT 47.68 51.439 55.356 54.444 ;
      RECT 0.7 0.986 55.356 54.158 ;
      RECT 0.7 0.7 19.776 3.705 ;
      RECT 41.904 0.7 55.356 3.705 ;
      POLYGON 32.544 55.144 32.544 55.088 32.388 55.088 32.388 54.444 32.544 54.444 32.544 54.158 34 54.158 34 54.444 38.32 54.444 38.32 54.158 39.776 54.158 39.776 54.444 40.448 54.444 40.448 54.158 41.904 54.158 41.904 54.444 42.576 54.444 42.576 54.158 44.032 54.158 44.032 54.444 46.224 54.444 46.224 54.158 47.68 54.158 47.68 54.444 55.356 54.444 55.356 0.7 41.904 0.7 41.904 0.986 40.448 0.986 40.448 0.7 39.776 0.7 39.776 0.986 38.32 0.986 38.32 0.7 36.128 0.7 36.128 0.986 34.672 0.986 34.672 0.7 34 0.7 34 0.986 32.544 0.986 32.544 0.7 31.872 0.7 31.872 0.986 30.416 0.986 30.416 0.7 29.744 0.7 29.744 0.986 28.288 0.986 28.288 0.7 28.132 0.7 28.132 0.191 28.134 0.191 28.134 0.081 28.074 0.081 28.074 0.191 28.076 0.191 28.076 0.7 27.616 0.7 27.616 0.986 26.16 0.986 26.16 0.7 25.7 0.7 25.7 0.191 25.702 0.191 25.702 0.081 25.642 0.081 25.642 0.191 25.644 0.191 25.644 0.7 25.488 0.7 25.488 0.986 24.032 0.986 24.032 0.7 23.36 0.7 23.36 0.986 21.904 0.986 21.904 0.7 21.444 0.7 21.444 0.108 21.232 0.108 21.232 0.164 21.388 0.164 21.388 0.7 21.232 0.7 21.232 0.986 19.776 0.986 19.776 0.7 0.7 0.7 0.7 54.444 15.52 54.444 15.52 54.158 16.976 54.158 16.976 54.444 25.856 54.444 25.856 54.158 27.312 54.158 27.312 54.444 32.332 54.444 32.332 55.144 ;
      RECT 0.106 26.676 0.166 26.943 ;
      POLYGON 55.95 21.471 55.95 21.361 55.948 21.361 55.948 21.167 55.95 21.167 55.95 21.057 55.89 21.057 55.89 21.167 55.892 21.167 55.892 21.361 55.89 21.361 55.89 21.471 ;
    LAYER M6 ;
      RECT 26.4 0.7 27.376 1.005 ;
      RECT 28.832 0.7 31.024 2.205 ;
      RECT 32.48 0.7 34.064 2.205 ;
      RECT 0.7 0.986 55.356 54.444 ;
      RECT 0.7 0.7 24.944 3.705 ;
      RECT 35.52 0.7 55.356 3.705 ;
    LAYER M3 ;
      RECT 55.051 44.336 55.356 45.008 ;
      RECT 55.051 41.904 55.356 42.88 ;
      RECT 55.051 39.776 55.356 40.448 ;
      RECT 55.051 37.04 55.356 38.32 ;
      RECT 55.051 34.912 55.356 35.584 ;
      RECT 55.051 32.784 55.356 33.456 ;
      RECT 0.7 32.176 1.005 32.848 ;
      RECT 55.051 30.048 55.356 31.328 ;
      RECT 0.7 30.048 1.005 30.72 ;
      RECT 0.7 27.92 1.005 28.592 ;
      RECT 55.051 27.312 55.356 28.592 ;
      RECT 55.051 21.84 55.356 22.512 ;
      RECT 55.051 19.712 55.356 20.384 ;
      RECT 0.7 24.272 2.205 26.464 ;
      RECT 53.851 23.968 55.356 25.856 ;
      RECT 0.7 20.928 2.205 22.816 ;
      RECT 0.7 46.464 55.356 54.444 ;
      RECT 0.7 34.304 55.07 46.464 ;
      RECT 0.986 19.472 55.07 34.304 ;
      RECT 0.986 18.256 55.07 21.261 ;
      RECT 0.7 16.467 3.705 19.472 ;
      RECT 0.7 0.7 55.356 18.256 ;
      POLYGON 55.356 54.444 55.356 46.464 55.07 46.464 55.07 45.008 55.356 45.008 55.356 44.336 55.07 44.336 55.07 42.88 55.356 42.88 55.356 41.904 55.07 41.904 55.07 40.448 55.356 40.448 55.356 39.776 55.07 39.776 55.07 38.32 55.356 38.32 55.356 37.04 55.07 37.04 55.07 35.584 55.356 35.584 55.356 34.912 55.07 34.912 55.07 33.456 55.356 33.456 55.356 32.784 55.07 32.784 55.07 31.328 55.356 31.328 55.356 30.048 55.07 30.048 55.07 28.592 55.356 28.592 55.356 27.312 55.07 27.312 55.07 25.856 55.356 25.856 55.356 23.968 55.07 23.968 55.07 22.512 55.356 22.512 55.356 21.84 55.07 21.84 55.07 20.384 55.356 20.384 55.356 19.712 55.07 19.712 55.07 18.256 55.356 18.256 55.356 0.7 0.7 0.7 0.7 19.472 0.986 19.472 0.986 20.928 0.7 20.928 0.7 22.816 0.986 22.816 0.986 24.272 0.7 24.272 0.7 26.464 0.986 26.464 0.986 26.86 0.191 26.86 0.191 26.858 0.081 26.858 0.081 26.918 0.191 26.918 0.191 26.916 0.986 26.916 0.986 27.92 0.7 27.92 0.7 28.592 0.986 28.592 0.986 30.048 0.7 30.048 0.7 30.72 0.986 30.72 0.986 32.176 0.7 32.176 0.7 32.848 0.986 32.848 0.986 34.304 0.7 34.304 0.7 54.444 ;
    LAYER M5 ;
      RECT 0.7 27.616 55.356 54.444 ;
      RECT 0.986 24.611 55.356 29.165 ;
      RECT 0.7 0.7 55.356 26.16 ;
      POLYGON 55.356 54.444 55.356 21.444 55.865 21.444 55.865 21.446 55.975 21.446 55.975 21.386 55.865 21.386 55.865 21.388 55.356 21.388 55.356 0.7 0.7 0.7 0.7 26.16 0.986 26.16 0.986 27.616 0.7 27.616 0.7 54.444 ;
      RECT 27.892 0.106 28.159 0.166 ;
      RECT 25.46 0.106 25.727 0.166 ;
    LAYER M8 ;
      RECT 0.7 53.444 0.9 54.444 ;
      RECT 55.156 53.444 55.356 54.444 ;
      RECT 0.7 0.7 0.9 1.7 ;
      RECT 55.156 0.7 55.356 1.7 ;
      RECT 4.7 51.439 51.356 54.444 ;
      RECT 0.7 1.7 55.356 53.444 ;
      RECT 4.7 0.7 51.356 3.705 ;
    LAYER M9 ;
      RECT 0.5 54.044 1.5 54.644 ;
      RECT 54.556 54.044 55.556 54.644 ;
      RECT 0.5 0.5 1.5 1.1 ;
      RECT 54.556 0.5 55.556 1.1 ;
      RECT 1.5 50.644 54.556 54.644 ;
      RECT 0.5 4.5 55.556 50.644 ;
      RECT 1.5 0.5 54.556 4.5 ;
    LAYER NWELL ;
      RECT 0.23 0.23 55.826 54.914 ;
    LAYER PO ;
      RECT 0.122 0.122 55.934 55.022 ;
    LAYER M1 ;
      RECT 0.6 0.6 55.456 54.544 ;
    LAYER M2 ;
      RECT 0.7 0.7 55.356 54.444 ;
    LAYER VIA3 ;
      RECT 0.111 26.863 0.161 26.913 ;
      RECT 55.895 21.087 55.945 21.137 ;
    LAYER VIA4 ;
      RECT 0.111 26.863 0.161 26.913 ;
      RECT 55.895 21.391 55.945 21.441 ;
      RECT 28.079 0.111 28.129 0.161 ;
      RECT 25.647 0.111 25.697 0.161 ;
    LAYER VIA5 ;
      RECT 28.079 0.111 28.129 0.161 ;
      RECT 25.647 0.111 25.697 0.161 ;
    LAYER M7 ;
      RECT 0.7 0.7 55.356 54.444 ;
    LAYER VIA8 ;
      RECT 54.266 53.354 54.396 53.484 ;
      RECT 54.016 53.354 54.146 53.484 ;
      RECT 53.766 53.354 53.896 53.484 ;
      RECT 53.516 53.354 53.646 53.484 ;
      RECT 2.41 53.354 2.54 53.484 ;
      RECT 2.16 53.354 2.29 53.484 ;
      RECT 1.91 53.354 2.04 53.484 ;
      RECT 1.66 53.354 1.79 53.484 ;
      RECT 54.266 1.66 54.396 1.79 ;
      RECT 54.016 1.66 54.146 1.79 ;
      RECT 53.766 1.66 53.896 1.79 ;
      RECT 53.516 1.66 53.646 1.79 ;
      RECT 2.41 1.66 2.54 1.79 ;
      RECT 2.16 1.66 2.29 1.79 ;
      RECT 1.91 1.66 2.04 1.79 ;
      RECT 1.66 1.66 1.79 1.79 ;
    LAYER MRDL ;
      RECT 2 2 54.056 53.144 ;
    LAYER OVERLAP ;
      POLYGON 0 0 0 55.144 56.056 55.144 56.056 0 ;
  END
END UART

END LIBRARY
